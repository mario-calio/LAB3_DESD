`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
gBARjbt2sG+aG4Anx+y0rKzF2Wd8e81IFJBsWFsXVGi3KxdrE9u/gOyyQSM2NjQI+jBc61yLelNf
YcTgu0NvLJs4vEEwWtZy1IfZLnvP83DlcPVVJK0YnXU2GXr4kBqtYMOkXtjtTJDoQHAY+RnvH39Y
typ2Kap1cY9uiKnMqK+gdhZxIKjpT/4ICJOi8TiGjkMLneYi0zy+Chm0VSQwA8rPO7ddXbjbr0+S
s7+JIcD+pV3heOvG7vHnTVbmb4miVgjT9WmUIDoodkIGVuavtfTxwPWlkm5SEBA3uO0B0c8wwRVA
Ps9byHhNhsggjRv1q2GOGAqToT/wiy0W3UYS7Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = "true"
`protect end_toolblock="lK7i8BiLYXJcsUUhiFTjcNrLKLCDf4VdoyV4twEGVI0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4128)
`protect data_block
JkuhdndhjqIA+liQHF1R86kXvR2J8m9t2Pitn7jKk7OuVgItMv/j6Xfst2KTKSorHwbzwCVVUwDs
roawsaxe5sfSUUhTnyz5lYRihHmwY1HSdI24S2E4E00f3OFmf9pv9BnV3xtCiQxO4jbfx3pZmFbK
ptdEwDMc2BEJDTyIubcdVqp4wu+51azrkkmZZcypxFfGbF8+Yi8hdcavbmm1MAv6Y0OCoFRe5Dke
dsoJf9peG8O9DB++LDnq6QIOIVknGFVReS0oqU3vZDKamJhq/xfggOIKo8yimXsD9qUZ4FgANkNH
XEPt7WKTjo9mzgQtW+D+KFvkUtTUh/WDfi04Gc93MYzoiiaiLYURHkXgbkadm2SVJo44n64/43Yu
8KX8J8KJhN6nIWWh91UYTRoiU2o6E2TGnJs/+WNAdEX7GLVswQRfLDD+vMtJrVcJSA2Cca68/TWD
2t28VigZOmXJVkAwY1h5KHMb96Ekl37C+TpcUtid3gRsDwSK0jdGYmRQo8myLhZt9bgnS/wAgn4y
tLbvY24S3OSL1eqInW48o8Tcug8Pvka2CV+VFS0mcGIY8GA9y3kxtpOMHqncN1HZx3c2reH5CT43
CurIUaq3v1oZC1sA9JrUtPnwng6DDPH2TgVSoF9+s/4b2h3o/i2/I03zdPc5wwSb3ApyXcUkUCw8
2ljKICGdCo8FEgk1YKPea8QJYk2a9Iffs5TqvNqBtm+okxtOGjLdrZ5PiQZw77gTLG8m5Y+RYhX+
NS0m2KUPEvwEtJGyuXRH4IqduDuV5eJ2Q9L36fNaE6+Juyi0v1Pr+IkhSKPZdf3pYQWDzujFWr5m
Pd7w7z0Z9eKQvqlHvp8sNfLVbfRQSba9fOExvwqe4WQWeM5RtwegTouKNerOTFHq8bc5qN7P+mbi
ZiUEcIEiya5OmjIX7Lsni84VeN1soo421ohLmRFNSH6W+ku/v/WOvt3AXXIjQ1cICuFATP/rXGIL
t0DUXZNGJX3xu2U1kdh5uIxlLojbaHP3MvDSUQ1b81YASJlwEqjDRVTKeye1qQ397xk4JRlVA4hZ
a2h1N1l28dXi2/wwgf/d5nsrXwLnavLpwdSps6loJbjEMdqTfNvDnMJzCNwaWGkIaoWAZvgPdFuR
zRs7BtmsaXr1PJzuFwbHOJ+xXFzGZ+bLgCSRL6HYyIprMELu2hO4bWpGKN9LPlN3fWPkGrXRE7sm
anGpPugqYHCO8fXswLrgkRq7HBREcuGRXoqZ5/BB1DZYM23iJz5DRKbOHaxUSNLIf59wy0qtUokx
hUzZNZ0dmdBdTXBIQDfrP/CdkS0Q0oJUh/FdvyY5GMMdem2+l51cwx7+xifmpPFL/Tk0ThH0KyXG
ckgqWUuHv/JhqLZfpglKNGjeQxJD7P9M40qNeQhiOJB4RRee4mVP3NahxYquCf/uCiI3mK2cmplQ
tUZpVt5tLA3vxEd/9KWq4uEFjnrNwZ6FmUqSaum6JDK0ruC34wKhyVUkp2Xwu15viXHNL1Zaisib
stWSNpMO7nS/6S9/KUD0ZjXu/3Tf7Dosg+lWy4AW74bKu3CgBlDbIMIQF3uPHCmbbv/7GsraXdDo
dFPQWFXG5EBO4RY01U2D4x3FJZzDbmzHJEpnKD9TSFYTF/vAHlqLsoaMRRQKEVaAeWPI8msUFazk
HFgMNwrKrczDQsHsgYYNlhPdBujHVTIQFP3j7/uBQaLyrOt4tjH5cve+U/GxE976mQpZv0QQ8Rv1
o7L1WRndHpT2StoPFVU1qB9qr7Sdi8yefI/tMs3YEmJeN8EprswtSYGtE84Z11j1BTNkOtp979OC
8CY+M6Xx071sKt0C8XIU9Ry1nXMnVdvAkIgjQo/tYWp+pDmTAHf+XBrW5uczfxMN7ItFL3an12MM
jAqiY5AbHg3JpiAdylGhYZGmYuEW2KFLBi6TSIWCqkW1d+RrdtY4NsFPzjjx5/X1N/YXiERBMcw5
YbbqJcC6pxGOH2P4s8VYgVSdKYGl3m391Q/UldR/0bbb6L+10t30YhP1Ocadl0YL1LUWIRPcSabv
qnE3RrhjBK7r9A7WdiikKiDQvCTRtgBLcbcMMf/4lIdKjXTPXfiXwyMJf6h7VGB5ovv9fXgGn3En
+prG76gw5bPixe8zd6FXuZ9hHosIQyxlT3vIRAYFFO71unUT1LovQ5zRwsvwF5Ji477Dyf9KGg5r
CVplzJN6kpb8Nd5bWD/7/q/beUI0YUgqRkGTEs0PF0Eg0xVMKeus7RZ+4MHoTepHMEaRILSaHw6h
XcYY0TBu159n5f1jLyCKo3WsH8b7IRGMqnGHYPTvCuMoQwLJJf0p+z4APMvsVWXSlcgqUJEtHxve
hM1SG/VSzKpxfb5e4rmT+CaH9VTAxntzQzlFaFD+MJWbySNVuokotni39abwxC1EEE47Fw/Qo+nd
s/xIcxaPtoHpdqoon2eHgORfotsNIeyBb3u9J7rhgWry9IVP3xbu6ow8DFeY+d0B2r2NmJtw/GmJ
DDVUkIqEqcqeTag0qY9/NhC9dU8sPjfRSMMaGb3OdAmy9pzV7I+AEb3AcyT0F7Lzb/vBPSJ6Mm4g
PGrp7IflztejMN7AAOI+QoG5SplcjxrYD5vGVjft61eh+JR5WPKcVbE057I6PiUHx56jwi+boMVd
w7RIKOd/8+47lNYlc99yvXnunCFRLI08+uUSEJ5f48+AGMpGLrj6BlOYxcD7hEwioCnqv50892r8
617qdweGi9AZmhwoLj9l9hf3+4CFSb9oaGKI6TP1k0D1ByxQ36BZw6QtB/n7KSADBXh3b5dEF1aJ
62MwCDy/xr4W6qvgaF4y5iy29z9TQGwr9mEjlXglb+TM5ecG2AgOwQaxj1VMCzSYezTET9RzVgr/
udJB7jbu2wKOFw9ogzmir0uZgVC6YCOHWf+rqQapw2jkQDiYzGmEf1Pee6jJq0EerI5WTuHLfYoo
BHHJb8J+q14fxHzNAJML6PcquHaLQBfDyJADFvYnGLizbwtKuCgHXJWtij6SpPgCfCrBJH2exRw8
LUllMufK2oM8UgDISsm7DelmSV04JjW+csYWUnrgqSRpJFCS/AxHSCd0o8UakjddWoupZmLvi3o6
MHFPtqS9rnQEtn8TeP8iODpP3ITP98CzCbucNmHYNLbk8+AEuVne0Q9dfei7T+1xj6H2v/vtWY6I
8rgdAGDeJHIuDb+zXzlgTDv+jkXjq4T4ERv9ZSv9GGXkJ86BVN3yewM+3Qa0ozqe12pwT3Od9cDG
9UuoCNOlv4gh4Fx9sofu1PoM3gmcDk43tOfKdhsjE2y/xXEcYsZP+BQrKHEBXj3qPA3v8s40Ridp
+vEkTexSmJfPekx96GWwaFCjAIZdqCRhMyxvHZBkgEBBUS99kgTDkQbenQJz9U8UD3yGDyxEqypR
cuIe6FhhZgN5qZg6fkQ51QuFD9h2lorVcAEkly1pV4yPHic9Lbhz0pCKmUU95g/rAglpRqdp8Q6Q
V/wGu5nL/++e25S8rbRdNSRB5fkcd5Zwu9XJ4j6gdQYSSbjerzVG4/Htt/NoDWTstETubVzaAopq
/X9fK1n1RwTP6NZMzJcZktJ5ijCdn9lD2dJXbtyAJSZVgEwNPZWGAHGjg5ClRbfyWb/kYpG0gSFa
Y78AIZ7lSiyjneRSTgVgLdb4Dv2HDEeuoNjoUWCLnKTxyvf1t/ZieksnCTqWIUnI2uxByMq9pLwN
0xJAMlJz4KPLkGq7cO0NYeC3yZEOfeu7cAEqFFBtCZCy2Y8xgh7Y5jzXMhYq/grsDVwjUR61Oqeh
3+3eawm6lV/hiyJlqMv27tZJrnrh81PPCdVXO5K2c2+ZwtCIBXNdYQY5tMquco6E8/DNz4xmB5Sx
Vh3MBb4VYYuzQpWFpp9XEfCjgA7FSP3Dq1sZR24wiPP6zN0g2m9mgeK4e0icCR9KlzitGpQn8pDF
n1X3LU1VIMP97ObfiQJk6fJHWhTN+gBjIeoWb3bwECOgrqbUJO9TEJjNuSLZUutViwqJLMSeYHgK
KwsGRwgWABTwRyXN9rcjyAWzl0V3qlZiSzyquW6awGaKdXz+ZfS6T+BGubWdgz8hesxGP95VrRB3
bZolMUfMByn8uW8LLUUtFoEVGDaXj6ML7zMNzBJjZ/tdw38L2ZhTJnWiO8rNxzJijlt2tt45z/kv
nW91nOWiqjFbQZ8cUU6bxuBOf6s/8ChHHaR7YUzLTjA/+55DiHxjLVAV5ik6Jv2BK7T/WsA9PEg6
GKXPOIrlXCwo4ANRN9F1xR75DuKocg6y/CQgxalfh189U+963lFf5PiBUC2xbFJuHtvwW7MiVsF4
lmJwAWdK8SLOjo0FW0XqVOqcp9+moT4YrU2WpXOcT8+GEsFb9M4E38S8AfVlEJxndIDOCeWaOVuz
9QTPPQ9NmINx3CInPE9qeiCNTvLaImTUepC0XK/q1W6NVzAMrYtKk61tlMPtV9vQAxB8R/58l3eb
lj3ITOLmczpVKKOvi4FDn2V9f2ry08RKD7gYAKNKIU3GMbHT00RqbRMJQJpMSQK7R6CQuVlSGWbM
R9DQb03bukrMuuNmKCS+wMQx70b9VX3QFtgip9aTBg/tSfmUl6wVGXkbNtSuehL5thA38Wx2w0JD
SN7apMExiSIkZwo+vaEtxtJpN33b+tsnuOtAWNSQsO+SJLHTX+sEjLe3zX1pJ0lGOyT8t9cRx9ra
8BT8alhE9ztJlsMhx9XALkXzaBn0ZwDHh+l1PTU6uVp3UjUEWrz+tjYmOsgV/eQXMYBnwF9PgFbK
qPNKy3QZFIhQzK/QjPYx6PCEggyVf8idSOmwXWgRGD/tjz8TEQcudU4WoAQ8Be6OARqXWF8XILjc
44lO1J18zeNnwgYnXbDdw83mpxVGWXhzB+XWnCGuGmtAvRGk3oTQacEGMDRDFEyflhmFVIEo9Hm0
IiJ8dg/3fjb1dnvRp3+spIR7wGCIJ4A0xK2XMhLDuHheVWfNf1ggljMHAweIWkENR987ofHXhzuD
l2KoyOcedQZ9tKsysYjKpHq2u1QwpJJCeQPS7H5fcZyn9fJeUynsULRaAa6OkgOdXse4JhuP/wgd
r172oggVK1SeXEzW9T3PTt2bsuy7Yc1teSMBHSwbQEqBDqwv7FB6iRd59xWRcBO/RcKWUWxvi5H+
u8n/i0HnsQnj6j9y/4RCrSGc20M5P3oryYP/nVhKvXZJvMwTru/FfKxVL/VQs0R0hvFU0hPdXhOD
QLPS2vee4sT18BOHMKWZBZxn5TALxju1zZy7MoNJPYwK4IXV1p7jX9sOIf8yHaH0Ia/NIkvkaZg2
jA0XZtnRHANDYopDnf+Os4ItFt12i9/ubfRWVZ74V2ixXVRONAYK+QWQG4NXQtJvcxnWg03eRKSZ
r5vYfcU8BG8OURvYvnaeEkQSMb0qId4Xg/CZMnI9LZC5Y+PJURxmsnBNg6uieGpP8JcDCCCqIgxa
HmtQHJIvqr9F3O7YUe1hx3kgxrB8bOvX
`protect end_protected
